** Profile: "SCHEMATIC1-Part1"  [ C:\USERS\ASUS\DESKTOP\H2\test-SCHEMATIC1-Part1.sim ] 

** Creating circuit file "test-SCHEMATIC1-Part1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\test-SCHEMATIC1.net" 


.END
