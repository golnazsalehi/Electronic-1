** Profile: "SCHEMATIC1-qesmat5"  [ c:\users\asus\desktop\elec\h1-SCHEMATIC1-qesmat5.sim ] 

** Creating circuit file "h1-SCHEMATIC1-qesmat5.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 0.001ms 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\h1-SCHEMATIC1.net" 


.END
