** Profile: "SCHEMATIC1-Real_part4"  [ c:\users\asus\desktop\h3\h3-schematic1-real_part4.sim ] 

** Creating circuit file "h3-schematic1-real_part4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 1k 30k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\h3-SCHEMATIC1.net" 


.END
