** Profile: "SCHEMATIC1-Part3"  [ c:\users\asus\desktop\h2\h2-SCHEMATIC1-Part3.sim ] 

** Creating circuit file "h2-SCHEMATIC1-Part3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1.5ms 0 0.0001ms 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\h2-SCHEMATIC1.net" 


.END
